`timescale 1ns/1ps
`include "../header_files/parameters.vh"

module stand_mode_controller_from_clean (
    input clk,      //100MHz clock signal
    input rstn,     //active-low
    input [`MODE_WIDTH-1:0] current_mode, // current mode
    output reg stand_mode_controller_from_clean_toggle // output toggle signal
);

reg turn_on_toggle_signal;
reg reset_timer_signal;
wire [`MAX_WIDTH-1:0] count_reg;
wire done;

countdown_timer from_clean_to_stand_timer_inst (
    .clk(clk),
    .rstn(rstn),
    .start(turn_on_toggle_signal),
    .load_value(`CLEAN_MODE_COUNTER_TIME),
    .reset_signal(reset_timer_signal),
    .count_reg(count_reg),
    .done(done)
);
reg started;
always @(posedge clk or negedge rstn) begin
    if (!rstn) begin
        stand_mode_controller_from_clean_toggle <= 1'b0;
        turn_on_toggle_signal <= 1'b0;
        reset_timer_signal <= 1'b1;
        started <= 1'b0;
    end else begin
        case (current_mode)
            `CLEAN_MODE: begin
                if (!done) begin
                    started <= 1'b1;
                end else if (done && !turn_on_toggle_signal) begin
                    turn_on_toggle_signal <= 1'b1;
                end else if (done && started) begin
                    stand_mode_controller_from_clean_toggle <= 1'b1;
                end
            end
            default: begin
                stand_mode_controller_from_clean_toggle <= 1'b0;
                turn_on_toggle_signal <= 1'b0;
                started <= 1'b0;
            end
        endcase
    end
end

endmodule //stand_mode_controller_from_clean