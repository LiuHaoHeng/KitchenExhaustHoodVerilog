`define OFF_MODE    8'b00000001
`define STAND_MODE  8'b00000010
`define CLEAN_MODE  8'b00000100
`define FIRST_MODE  8'b00001000 
`define SECOND_MODE 8'b00010000 
`define THIRD_MODE  8'b00100000  
`define SET_MODE    8'b01000000
`define PRE_MODE    8'b10000000

`define MODE_WIDTH 8

`define MAX_WIDTH 32
`define COUNTER_1SEC 100000000

`define OFF_MODE_NORMAL_COUNT_TIME 300000000
`define OFF_MODE_GESTURE_COUNTER_TIME 5

`define CLEAN_MODE_COUNTER_TIME 10
`define THIRD_MODE_COUNTER_TIME 7

`define OUTPUT_WIDTH 8

`define MAX_GESTURE_TIME 32'd7
`define DEFAULT_GESTURE_TIME 32'd5
`define MIN_GESTURE_TIME 32'd2
    
`define MAX_CLEAN_REMIND_TIME 32'd108000
`define DEFAULT_CLEAN_REMIND_TIME 32'd36000
`define MIN_CLEAN_REMIND_TIME 32'd10